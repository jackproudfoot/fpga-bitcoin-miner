module reg640(q, d, clk, en, clr);
	input [639:0] d; 
	input clk, en, clr;
	output [639:0] q;

	dffe_ref flipFlop0(q[0], d[0], clk, en, clr);
	dffe_ref flipFlop1(q[1], d[1], clk, en, clr);
	dffe_ref flipFlop2(q[2], d[2], clk, en, clr);
	dffe_ref flipFlop3(q[3], d[3], clk, en, clr);
	dffe_ref flipFlop4(q[4], d[4], clk, en, clr);
	dffe_ref flipFlop5(q[5], d[5], clk, en, clr);
	dffe_ref flipFlop6(q[6], d[6], clk, en, clr);
	dffe_ref flipFlop7(q[7], d[7], clk, en, clr);
	dffe_ref flipFlop8(q[8], d[8], clk, en, clr);
	dffe_ref flipFlop9(q[9], d[9], clk, en, clr);
	dffe_ref flipFlop10(q[10], d[10], clk, en, clr);
	dffe_ref flipFlop11(q[11], d[11], clk, en, clr);
	dffe_ref flipFlop12(q[12], d[12], clk, en, clr);
	dffe_ref flipFlop13(q[13], d[13], clk, en, clr);
	dffe_ref flipFlop14(q[14], d[14], clk, en, clr);
	dffe_ref flipFlop15(q[15], d[15], clk, en, clr);
	dffe_ref flipFlop16(q[16], d[16], clk, en, clr);
	dffe_ref flipFlop17(q[17], d[17], clk, en, clr);
	dffe_ref flipFlop18(q[18], d[18], clk, en, clr);
	dffe_ref flipFlop19(q[19], d[19], clk, en, clr);
	dffe_ref flipFlop20(q[20], d[20], clk, en, clr);
	dffe_ref flipFlop21(q[21], d[21], clk, en, clr);
	dffe_ref flipFlop22(q[22], d[22], clk, en, clr);
	dffe_ref flipFlop23(q[23], d[23], clk, en, clr);
	dffe_ref flipFlop24(q[24], d[24], clk, en, clr);
	dffe_ref flipFlop25(q[25], d[25], clk, en, clr);
	dffe_ref flipFlop26(q[26], d[26], clk, en, clr);
	dffe_ref flipFlop27(q[27], d[27], clk, en, clr);
	dffe_ref flipFlop28(q[28], d[28], clk, en, clr);
	dffe_ref flipFlop29(q[29], d[29], clk, en, clr);
	dffe_ref flipFlop30(q[30], d[30], clk, en, clr);
	dffe_ref flipFlop31(q[31], d[31], clk, en, clr);
	dffe_ref flipFlop32(q[32], d[32], clk, en, clr);
	dffe_ref flipFlop33(q[33], d[33], clk, en, clr);
	dffe_ref flipFlop34(q[34], d[34], clk, en, clr);
	dffe_ref flipFlop35(q[35], d[35], clk, en, clr);
	dffe_ref flipFlop36(q[36], d[36], clk, en, clr);
	dffe_ref flipFlop37(q[37], d[37], clk, en, clr);
	dffe_ref flipFlop38(q[38], d[38], clk, en, clr);
	dffe_ref flipFlop39(q[39], d[39], clk, en, clr);
	dffe_ref flipFlop40(q[40], d[40], clk, en, clr);
	dffe_ref flipFlop41(q[41], d[41], clk, en, clr);
	dffe_ref flipFlop42(q[42], d[42], clk, en, clr);
	dffe_ref flipFlop43(q[43], d[43], clk, en, clr);
	dffe_ref flipFlop44(q[44], d[44], clk, en, clr);
	dffe_ref flipFlop45(q[45], d[45], clk, en, clr);
	dffe_ref flipFlop46(q[46], d[46], clk, en, clr);
	dffe_ref flipFlop47(q[47], d[47], clk, en, clr);
	dffe_ref flipFlop48(q[48], d[48], clk, en, clr);
	dffe_ref flipFlop49(q[49], d[49], clk, en, clr);
	dffe_ref flipFlop50(q[50], d[50], clk, en, clr);
	dffe_ref flipFlop51(q[51], d[51], clk, en, clr);
	dffe_ref flipFlop52(q[52], d[52], clk, en, clr);
	dffe_ref flipFlop53(q[53], d[53], clk, en, clr);
	dffe_ref flipFlop54(q[54], d[54], clk, en, clr);
	dffe_ref flipFlop55(q[55], d[55], clk, en, clr);
	dffe_ref flipFlop56(q[56], d[56], clk, en, clr);
	dffe_ref flipFlop57(q[57], d[57], clk, en, clr);
	dffe_ref flipFlop58(q[58], d[58], clk, en, clr);
	dffe_ref flipFlop59(q[59], d[59], clk, en, clr);
	dffe_ref flipFlop60(q[60], d[60], clk, en, clr);
	dffe_ref flipFlop61(q[61], d[61], clk, en, clr);
	dffe_ref flipFlop62(q[62], d[62], clk, en, clr);
	dffe_ref flipFlop63(q[63], d[63], clk, en, clr);
	dffe_ref flipFlop64(q[64], d[64], clk, en, clr);
	dffe_ref flipFlop65(q[65], d[65], clk, en, clr);
	dffe_ref flipFlop66(q[66], d[66], clk, en, clr);
	dffe_ref flipFlop67(q[67], d[67], clk, en, clr);
	dffe_ref flipFlop68(q[68], d[68], clk, en, clr);
	dffe_ref flipFlop69(q[69], d[69], clk, en, clr);
	dffe_ref flipFlop70(q[70], d[70], clk, en, clr);
	dffe_ref flipFlop71(q[71], d[71], clk, en, clr);
	dffe_ref flipFlop72(q[72], d[72], clk, en, clr);
	dffe_ref flipFlop73(q[73], d[73], clk, en, clr);
	dffe_ref flipFlop74(q[74], d[74], clk, en, clr);
	dffe_ref flipFlop75(q[75], d[75], clk, en, clr);
	dffe_ref flipFlop76(q[76], d[76], clk, en, clr);
	dffe_ref flipFlop77(q[77], d[77], clk, en, clr);
	dffe_ref flipFlop78(q[78], d[78], clk, en, clr);
	dffe_ref flipFlop79(q[79], d[79], clk, en, clr);
	dffe_ref flipFlop80(q[80], d[80], clk, en, clr);
	dffe_ref flipFlop81(q[81], d[81], clk, en, clr);
	dffe_ref flipFlop82(q[82], d[82], clk, en, clr);
	dffe_ref flipFlop83(q[83], d[83], clk, en, clr);
	dffe_ref flipFlop84(q[84], d[84], clk, en, clr);
	dffe_ref flipFlop85(q[85], d[85], clk, en, clr);
	dffe_ref flipFlop86(q[86], d[86], clk, en, clr);
	dffe_ref flipFlop87(q[87], d[87], clk, en, clr);
	dffe_ref flipFlop88(q[88], d[88], clk, en, clr);
	dffe_ref flipFlop89(q[89], d[89], clk, en, clr);
	dffe_ref flipFlop90(q[90], d[90], clk, en, clr);
	dffe_ref flipFlop91(q[91], d[91], clk, en, clr);
	dffe_ref flipFlop92(q[92], d[92], clk, en, clr);
	dffe_ref flipFlop93(q[93], d[93], clk, en, clr);
	dffe_ref flipFlop94(q[94], d[94], clk, en, clr);
	dffe_ref flipFlop95(q[95], d[95], clk, en, clr);
	dffe_ref flipFlop96(q[96], d[96], clk, en, clr);
	dffe_ref flipFlop97(q[97], d[97], clk, en, clr);
	dffe_ref flipFlop98(q[98], d[98], clk, en, clr);
	dffe_ref flipFlop99(q[99], d[99], clk, en, clr);
	dffe_ref flipFlop100(q[100], d[100], clk, en, clr);
	dffe_ref flipFlop101(q[101], d[101], clk, en, clr);
	dffe_ref flipFlop102(q[102], d[102], clk, en, clr);
	dffe_ref flipFlop103(q[103], d[103], clk, en, clr);
	dffe_ref flipFlop104(q[104], d[104], clk, en, clr);
	dffe_ref flipFlop105(q[105], d[105], clk, en, clr);
	dffe_ref flipFlop106(q[106], d[106], clk, en, clr);
	dffe_ref flipFlop107(q[107], d[107], clk, en, clr);
	dffe_ref flipFlop108(q[108], d[108], clk, en, clr);
	dffe_ref flipFlop109(q[109], d[109], clk, en, clr);
	dffe_ref flipFlop110(q[110], d[110], clk, en, clr);
	dffe_ref flipFlop111(q[111], d[111], clk, en, clr);
	dffe_ref flipFlop112(q[112], d[112], clk, en, clr);
	dffe_ref flipFlop113(q[113], d[113], clk, en, clr);
	dffe_ref flipFlop114(q[114], d[114], clk, en, clr);
	dffe_ref flipFlop115(q[115], d[115], clk, en, clr);
	dffe_ref flipFlop116(q[116], d[116], clk, en, clr);
	dffe_ref flipFlop117(q[117], d[117], clk, en, clr);
	dffe_ref flipFlop118(q[118], d[118], clk, en, clr);
	dffe_ref flipFlop119(q[119], d[119], clk, en, clr);
	dffe_ref flipFlop120(q[120], d[120], clk, en, clr);
	dffe_ref flipFlop121(q[121], d[121], clk, en, clr);
	dffe_ref flipFlop122(q[122], d[122], clk, en, clr);
	dffe_ref flipFlop123(q[123], d[123], clk, en, clr);
	dffe_ref flipFlop124(q[124], d[124], clk, en, clr);
	dffe_ref flipFlop125(q[125], d[125], clk, en, clr);
	dffe_ref flipFlop126(q[126], d[126], clk, en, clr);
	dffe_ref flipFlop127(q[127], d[127], clk, en, clr);
	dffe_ref flipFlop128(q[128], d[128], clk, en, clr);
	dffe_ref flipFlop129(q[129], d[129], clk, en, clr);
	dffe_ref flipFlop130(q[130], d[130], clk, en, clr);
	dffe_ref flipFlop131(q[131], d[131], clk, en, clr);
	dffe_ref flipFlop132(q[132], d[132], clk, en, clr);
	dffe_ref flipFlop133(q[133], d[133], clk, en, clr);
	dffe_ref flipFlop134(q[134], d[134], clk, en, clr);
	dffe_ref flipFlop135(q[135], d[135], clk, en, clr);
	dffe_ref flipFlop136(q[136], d[136], clk, en, clr);
	dffe_ref flipFlop137(q[137], d[137], clk, en, clr);
	dffe_ref flipFlop138(q[138], d[138], clk, en, clr);
	dffe_ref flipFlop139(q[139], d[139], clk, en, clr);
	dffe_ref flipFlop140(q[140], d[140], clk, en, clr);
	dffe_ref flipFlop141(q[141], d[141], clk, en, clr);
	dffe_ref flipFlop142(q[142], d[142], clk, en, clr);
	dffe_ref flipFlop143(q[143], d[143], clk, en, clr);
	dffe_ref flipFlop144(q[144], d[144], clk, en, clr);
	dffe_ref flipFlop145(q[145], d[145], clk, en, clr);
	dffe_ref flipFlop146(q[146], d[146], clk, en, clr);
	dffe_ref flipFlop147(q[147], d[147], clk, en, clr);
	dffe_ref flipFlop148(q[148], d[148], clk, en, clr);
	dffe_ref flipFlop149(q[149], d[149], clk, en, clr);
	dffe_ref flipFlop150(q[150], d[150], clk, en, clr);
	dffe_ref flipFlop151(q[151], d[151], clk, en, clr);
	dffe_ref flipFlop152(q[152], d[152], clk, en, clr);
	dffe_ref flipFlop153(q[153], d[153], clk, en, clr);
	dffe_ref flipFlop154(q[154], d[154], clk, en, clr);
	dffe_ref flipFlop155(q[155], d[155], clk, en, clr);
	dffe_ref flipFlop156(q[156], d[156], clk, en, clr);
	dffe_ref flipFlop157(q[157], d[157], clk, en, clr);
	dffe_ref flipFlop158(q[158], d[158], clk, en, clr);
	dffe_ref flipFlop159(q[159], d[159], clk, en, clr);
	dffe_ref flipFlop160(q[160], d[160], clk, en, clr);
	dffe_ref flipFlop161(q[161], d[161], clk, en, clr);
	dffe_ref flipFlop162(q[162], d[162], clk, en, clr);
	dffe_ref flipFlop163(q[163], d[163], clk, en, clr);
	dffe_ref flipFlop164(q[164], d[164], clk, en, clr);
	dffe_ref flipFlop165(q[165], d[165], clk, en, clr);
	dffe_ref flipFlop166(q[166], d[166], clk, en, clr);
	dffe_ref flipFlop167(q[167], d[167], clk, en, clr);
	dffe_ref flipFlop168(q[168], d[168], clk, en, clr);
	dffe_ref flipFlop169(q[169], d[169], clk, en, clr);
	dffe_ref flipFlop170(q[170], d[170], clk, en, clr);
	dffe_ref flipFlop171(q[171], d[171], clk, en, clr);
	dffe_ref flipFlop172(q[172], d[172], clk, en, clr);
	dffe_ref flipFlop173(q[173], d[173], clk, en, clr);
	dffe_ref flipFlop174(q[174], d[174], clk, en, clr);
	dffe_ref flipFlop175(q[175], d[175], clk, en, clr);
	dffe_ref flipFlop176(q[176], d[176], clk, en, clr);
	dffe_ref flipFlop177(q[177], d[177], clk, en, clr);
	dffe_ref flipFlop178(q[178], d[178], clk, en, clr);
	dffe_ref flipFlop179(q[179], d[179], clk, en, clr);
	dffe_ref flipFlop180(q[180], d[180], clk, en, clr);
	dffe_ref flipFlop181(q[181], d[181], clk, en, clr);
	dffe_ref flipFlop182(q[182], d[182], clk, en, clr);
	dffe_ref flipFlop183(q[183], d[183], clk, en, clr);
	dffe_ref flipFlop184(q[184], d[184], clk, en, clr);
	dffe_ref flipFlop185(q[185], d[185], clk, en, clr);
	dffe_ref flipFlop186(q[186], d[186], clk, en, clr);
	dffe_ref flipFlop187(q[187], d[187], clk, en, clr);
	dffe_ref flipFlop188(q[188], d[188], clk, en, clr);
	dffe_ref flipFlop189(q[189], d[189], clk, en, clr);
	dffe_ref flipFlop190(q[190], d[190], clk, en, clr);
	dffe_ref flipFlop191(q[191], d[191], clk, en, clr);
	dffe_ref flipFlop192(q[192], d[192], clk, en, clr);
	dffe_ref flipFlop193(q[193], d[193], clk, en, clr);
	dffe_ref flipFlop194(q[194], d[194], clk, en, clr);
	dffe_ref flipFlop195(q[195], d[195], clk, en, clr);
	dffe_ref flipFlop196(q[196], d[196], clk, en, clr);
	dffe_ref flipFlop197(q[197], d[197], clk, en, clr);
	dffe_ref flipFlop198(q[198], d[198], clk, en, clr);
	dffe_ref flipFlop199(q[199], d[199], clk, en, clr);
	dffe_ref flipFlop200(q[200], d[200], clk, en, clr);
	dffe_ref flipFlop201(q[201], d[201], clk, en, clr);
	dffe_ref flipFlop202(q[202], d[202], clk, en, clr);
	dffe_ref flipFlop203(q[203], d[203], clk, en, clr);
	dffe_ref flipFlop204(q[204], d[204], clk, en, clr);
	dffe_ref flipFlop205(q[205], d[205], clk, en, clr);
	dffe_ref flipFlop206(q[206], d[206], clk, en, clr);
	dffe_ref flipFlop207(q[207], d[207], clk, en, clr);
	dffe_ref flipFlop208(q[208], d[208], clk, en, clr);
	dffe_ref flipFlop209(q[209], d[209], clk, en, clr);
	dffe_ref flipFlop210(q[210], d[210], clk, en, clr);
	dffe_ref flipFlop211(q[211], d[211], clk, en, clr);
	dffe_ref flipFlop212(q[212], d[212], clk, en, clr);
	dffe_ref flipFlop213(q[213], d[213], clk, en, clr);
	dffe_ref flipFlop214(q[214], d[214], clk, en, clr);
	dffe_ref flipFlop215(q[215], d[215], clk, en, clr);
	dffe_ref flipFlop216(q[216], d[216], clk, en, clr);
	dffe_ref flipFlop217(q[217], d[217], clk, en, clr);
	dffe_ref flipFlop218(q[218], d[218], clk, en, clr);
	dffe_ref flipFlop219(q[219], d[219], clk, en, clr);
	dffe_ref flipFlop220(q[220], d[220], clk, en, clr);
	dffe_ref flipFlop221(q[221], d[221], clk, en, clr);
	dffe_ref flipFlop222(q[222], d[222], clk, en, clr);
	dffe_ref flipFlop223(q[223], d[223], clk, en, clr);
	dffe_ref flipFlop224(q[224], d[224], clk, en, clr);
	dffe_ref flipFlop225(q[225], d[225], clk, en, clr);
	dffe_ref flipFlop226(q[226], d[226], clk, en, clr);
	dffe_ref flipFlop227(q[227], d[227], clk, en, clr);
	dffe_ref flipFlop228(q[228], d[228], clk, en, clr);
	dffe_ref flipFlop229(q[229], d[229], clk, en, clr);
	dffe_ref flipFlop230(q[230], d[230], clk, en, clr);
	dffe_ref flipFlop231(q[231], d[231], clk, en, clr);
	dffe_ref flipFlop232(q[232], d[232], clk, en, clr);
	dffe_ref flipFlop233(q[233], d[233], clk, en, clr);
	dffe_ref flipFlop234(q[234], d[234], clk, en, clr);
	dffe_ref flipFlop235(q[235], d[235], clk, en, clr);
	dffe_ref flipFlop236(q[236], d[236], clk, en, clr);
	dffe_ref flipFlop237(q[237], d[237], clk, en, clr);
	dffe_ref flipFlop238(q[238], d[238], clk, en, clr);
	dffe_ref flipFlop239(q[239], d[239], clk, en, clr);
	dffe_ref flipFlop240(q[240], d[240], clk, en, clr);
	dffe_ref flipFlop241(q[241], d[241], clk, en, clr);
	dffe_ref flipFlop242(q[242], d[242], clk, en, clr);
	dffe_ref flipFlop243(q[243], d[243], clk, en, clr);
	dffe_ref flipFlop244(q[244], d[244], clk, en, clr);
	dffe_ref flipFlop245(q[245], d[245], clk, en, clr);
	dffe_ref flipFlop246(q[246], d[246], clk, en, clr);
	dffe_ref flipFlop247(q[247], d[247], clk, en, clr);
	dffe_ref flipFlop248(q[248], d[248], clk, en, clr);
	dffe_ref flipFlop249(q[249], d[249], clk, en, clr);
	dffe_ref flipFlop250(q[250], d[250], clk, en, clr);
	dffe_ref flipFlop251(q[251], d[251], clk, en, clr);
	dffe_ref flipFlop252(q[252], d[252], clk, en, clr);
	dffe_ref flipFlop253(q[253], d[253], clk, en, clr);
	dffe_ref flipFlop254(q[254], d[254], clk, en, clr);
	dffe_ref flipFlop255(q[255], d[255], clk, en, clr);
	dffe_ref flipFlop256(q[256], d[256], clk, en, clr);
	dffe_ref flipFlop257(q[257], d[257], clk, en, clr);
	dffe_ref flipFlop258(q[258], d[258], clk, en, clr);
	dffe_ref flipFlop259(q[259], d[259], clk, en, clr);
	dffe_ref flipFlop260(q[260], d[260], clk, en, clr);
	dffe_ref flipFlop261(q[261], d[261], clk, en, clr);
	dffe_ref flipFlop262(q[262], d[262], clk, en, clr);
	dffe_ref flipFlop263(q[263], d[263], clk, en, clr);
	dffe_ref flipFlop264(q[264], d[264], clk, en, clr);
	dffe_ref flipFlop265(q[265], d[265], clk, en, clr);
	dffe_ref flipFlop266(q[266], d[266], clk, en, clr);
	dffe_ref flipFlop267(q[267], d[267], clk, en, clr);
	dffe_ref flipFlop268(q[268], d[268], clk, en, clr);
	dffe_ref flipFlop269(q[269], d[269], clk, en, clr);
	dffe_ref flipFlop270(q[270], d[270], clk, en, clr);
	dffe_ref flipFlop271(q[271], d[271], clk, en, clr);
	dffe_ref flipFlop272(q[272], d[272], clk, en, clr);
	dffe_ref flipFlop273(q[273], d[273], clk, en, clr);
	dffe_ref flipFlop274(q[274], d[274], clk, en, clr);
	dffe_ref flipFlop275(q[275], d[275], clk, en, clr);
	dffe_ref flipFlop276(q[276], d[276], clk, en, clr);
	dffe_ref flipFlop277(q[277], d[277], clk, en, clr);
	dffe_ref flipFlop278(q[278], d[278], clk, en, clr);
	dffe_ref flipFlop279(q[279], d[279], clk, en, clr);
	dffe_ref flipFlop280(q[280], d[280], clk, en, clr);
	dffe_ref flipFlop281(q[281], d[281], clk, en, clr);
	dffe_ref flipFlop282(q[282], d[282], clk, en, clr);
	dffe_ref flipFlop283(q[283], d[283], clk, en, clr);
	dffe_ref flipFlop284(q[284], d[284], clk, en, clr);
	dffe_ref flipFlop285(q[285], d[285], clk, en, clr);
	dffe_ref flipFlop286(q[286], d[286], clk, en, clr);
	dffe_ref flipFlop287(q[287], d[287], clk, en, clr);
	dffe_ref flipFlop288(q[288], d[288], clk, en, clr);
	dffe_ref flipFlop289(q[289], d[289], clk, en, clr);
	dffe_ref flipFlop290(q[290], d[290], clk, en, clr);
	dffe_ref flipFlop291(q[291], d[291], clk, en, clr);
	dffe_ref flipFlop292(q[292], d[292], clk, en, clr);
	dffe_ref flipFlop293(q[293], d[293], clk, en, clr);
	dffe_ref flipFlop294(q[294], d[294], clk, en, clr);
	dffe_ref flipFlop295(q[295], d[295], clk, en, clr);
	dffe_ref flipFlop296(q[296], d[296], clk, en, clr);
	dffe_ref flipFlop297(q[297], d[297], clk, en, clr);
	dffe_ref flipFlop298(q[298], d[298], clk, en, clr);
	dffe_ref flipFlop299(q[299], d[299], clk, en, clr);
	dffe_ref flipFlop300(q[300], d[300], clk, en, clr);
	dffe_ref flipFlop301(q[301], d[301], clk, en, clr);
	dffe_ref flipFlop302(q[302], d[302], clk, en, clr);
	dffe_ref flipFlop303(q[303], d[303], clk, en, clr);
	dffe_ref flipFlop304(q[304], d[304], clk, en, clr);
	dffe_ref flipFlop305(q[305], d[305], clk, en, clr);
	dffe_ref flipFlop306(q[306], d[306], clk, en, clr);
	dffe_ref flipFlop307(q[307], d[307], clk, en, clr);
	dffe_ref flipFlop308(q[308], d[308], clk, en, clr);
	dffe_ref flipFlop309(q[309], d[309], clk, en, clr);
	dffe_ref flipFlop310(q[310], d[310], clk, en, clr);
	dffe_ref flipFlop311(q[311], d[311], clk, en, clr);
	dffe_ref flipFlop312(q[312], d[312], clk, en, clr);
	dffe_ref flipFlop313(q[313], d[313], clk, en, clr);
	dffe_ref flipFlop314(q[314], d[314], clk, en, clr);
	dffe_ref flipFlop315(q[315], d[315], clk, en, clr);
	dffe_ref flipFlop316(q[316], d[316], clk, en, clr);
	dffe_ref flipFlop317(q[317], d[317], clk, en, clr);
	dffe_ref flipFlop318(q[318], d[318], clk, en, clr);
	dffe_ref flipFlop319(q[319], d[319], clk, en, clr);
	dffe_ref flipFlop320(q[320], d[320], clk, en, clr);
	dffe_ref flipFlop321(q[321], d[321], clk, en, clr);
	dffe_ref flipFlop322(q[322], d[322], clk, en, clr);
	dffe_ref flipFlop323(q[323], d[323], clk, en, clr);
	dffe_ref flipFlop324(q[324], d[324], clk, en, clr);
	dffe_ref flipFlop325(q[325], d[325], clk, en, clr);
	dffe_ref flipFlop326(q[326], d[326], clk, en, clr);
	dffe_ref flipFlop327(q[327], d[327], clk, en, clr);
	dffe_ref flipFlop328(q[328], d[328], clk, en, clr);
	dffe_ref flipFlop329(q[329], d[329], clk, en, clr);
	dffe_ref flipFlop330(q[330], d[330], clk, en, clr);
	dffe_ref flipFlop331(q[331], d[331], clk, en, clr);
	dffe_ref flipFlop332(q[332], d[332], clk, en, clr);
	dffe_ref flipFlop333(q[333], d[333], clk, en, clr);
	dffe_ref flipFlop334(q[334], d[334], clk, en, clr);
	dffe_ref flipFlop335(q[335], d[335], clk, en, clr);
	dffe_ref flipFlop336(q[336], d[336], clk, en, clr);
	dffe_ref flipFlop337(q[337], d[337], clk, en, clr);
	dffe_ref flipFlop338(q[338], d[338], clk, en, clr);
	dffe_ref flipFlop339(q[339], d[339], clk, en, clr);
	dffe_ref flipFlop340(q[340], d[340], clk, en, clr);
	dffe_ref flipFlop341(q[341], d[341], clk, en, clr);
	dffe_ref flipFlop342(q[342], d[342], clk, en, clr);
	dffe_ref flipFlop343(q[343], d[343], clk, en, clr);
	dffe_ref flipFlop344(q[344], d[344], clk, en, clr);
	dffe_ref flipFlop345(q[345], d[345], clk, en, clr);
	dffe_ref flipFlop346(q[346], d[346], clk, en, clr);
	dffe_ref flipFlop347(q[347], d[347], clk, en, clr);
	dffe_ref flipFlop348(q[348], d[348], clk, en, clr);
	dffe_ref flipFlop349(q[349], d[349], clk, en, clr);
	dffe_ref flipFlop350(q[350], d[350], clk, en, clr);
	dffe_ref flipFlop351(q[351], d[351], clk, en, clr);
	dffe_ref flipFlop352(q[352], d[352], clk, en, clr);
	dffe_ref flipFlop353(q[353], d[353], clk, en, clr);
	dffe_ref flipFlop354(q[354], d[354], clk, en, clr);
	dffe_ref flipFlop355(q[355], d[355], clk, en, clr);
	dffe_ref flipFlop356(q[356], d[356], clk, en, clr);
	dffe_ref flipFlop357(q[357], d[357], clk, en, clr);
	dffe_ref flipFlop358(q[358], d[358], clk, en, clr);
	dffe_ref flipFlop359(q[359], d[359], clk, en, clr);
	dffe_ref flipFlop360(q[360], d[360], clk, en, clr);
	dffe_ref flipFlop361(q[361], d[361], clk, en, clr);
	dffe_ref flipFlop362(q[362], d[362], clk, en, clr);
	dffe_ref flipFlop363(q[363], d[363], clk, en, clr);
	dffe_ref flipFlop364(q[364], d[364], clk, en, clr);
	dffe_ref flipFlop365(q[365], d[365], clk, en, clr);
	dffe_ref flipFlop366(q[366], d[366], clk, en, clr);
	dffe_ref flipFlop367(q[367], d[367], clk, en, clr);
	dffe_ref flipFlop368(q[368], d[368], clk, en, clr);
	dffe_ref flipFlop369(q[369], d[369], clk, en, clr);
	dffe_ref flipFlop370(q[370], d[370], clk, en, clr);
	dffe_ref flipFlop371(q[371], d[371], clk, en, clr);
	dffe_ref flipFlop372(q[372], d[372], clk, en, clr);
	dffe_ref flipFlop373(q[373], d[373], clk, en, clr);
	dffe_ref flipFlop374(q[374], d[374], clk, en, clr);
	dffe_ref flipFlop375(q[375], d[375], clk, en, clr);
	dffe_ref flipFlop376(q[376], d[376], clk, en, clr);
	dffe_ref flipFlop377(q[377], d[377], clk, en, clr);
	dffe_ref flipFlop378(q[378], d[378], clk, en, clr);
	dffe_ref flipFlop379(q[379], d[379], clk, en, clr);
	dffe_ref flipFlop380(q[380], d[380], clk, en, clr);
	dffe_ref flipFlop381(q[381], d[381], clk, en, clr);
	dffe_ref flipFlop382(q[382], d[382], clk, en, clr);
	dffe_ref flipFlop383(q[383], d[383], clk, en, clr);
	dffe_ref flipFlop384(q[384], d[384], clk, en, clr);
	dffe_ref flipFlop385(q[385], d[385], clk, en, clr);
	dffe_ref flipFlop386(q[386], d[386], clk, en, clr);
	dffe_ref flipFlop387(q[387], d[387], clk, en, clr);
	dffe_ref flipFlop388(q[388], d[388], clk, en, clr);
	dffe_ref flipFlop389(q[389], d[389], clk, en, clr);
	dffe_ref flipFlop390(q[390], d[390], clk, en, clr);
	dffe_ref flipFlop391(q[391], d[391], clk, en, clr);
	dffe_ref flipFlop392(q[392], d[392], clk, en, clr);
	dffe_ref flipFlop393(q[393], d[393], clk, en, clr);
	dffe_ref flipFlop394(q[394], d[394], clk, en, clr);
	dffe_ref flipFlop395(q[395], d[395], clk, en, clr);
	dffe_ref flipFlop396(q[396], d[396], clk, en, clr);
	dffe_ref flipFlop397(q[397], d[397], clk, en, clr);
	dffe_ref flipFlop398(q[398], d[398], clk, en, clr);
	dffe_ref flipFlop399(q[399], d[399], clk, en, clr);
	dffe_ref flipFlop400(q[400], d[400], clk, en, clr);
	dffe_ref flipFlop401(q[401], d[401], clk, en, clr);
	dffe_ref flipFlop402(q[402], d[402], clk, en, clr);
	dffe_ref flipFlop403(q[403], d[403], clk, en, clr);
	dffe_ref flipFlop404(q[404], d[404], clk, en, clr);
	dffe_ref flipFlop405(q[405], d[405], clk, en, clr);
	dffe_ref flipFlop406(q[406], d[406], clk, en, clr);
	dffe_ref flipFlop407(q[407], d[407], clk, en, clr);
	dffe_ref flipFlop408(q[408], d[408], clk, en, clr);
	dffe_ref flipFlop409(q[409], d[409], clk, en, clr);
	dffe_ref flipFlop410(q[410], d[410], clk, en, clr);
	dffe_ref flipFlop411(q[411], d[411], clk, en, clr);
	dffe_ref flipFlop412(q[412], d[412], clk, en, clr);
	dffe_ref flipFlop413(q[413], d[413], clk, en, clr);
	dffe_ref flipFlop414(q[414], d[414], clk, en, clr);
	dffe_ref flipFlop415(q[415], d[415], clk, en, clr);
	dffe_ref flipFlop416(q[416], d[416], clk, en, clr);
	dffe_ref flipFlop417(q[417], d[417], clk, en, clr);
	dffe_ref flipFlop418(q[418], d[418], clk, en, clr);
	dffe_ref flipFlop419(q[419], d[419], clk, en, clr);
	dffe_ref flipFlop420(q[420], d[420], clk, en, clr);
	dffe_ref flipFlop421(q[421], d[421], clk, en, clr);
	dffe_ref flipFlop422(q[422], d[422], clk, en, clr);
	dffe_ref flipFlop423(q[423], d[423], clk, en, clr);
	dffe_ref flipFlop424(q[424], d[424], clk, en, clr);
	dffe_ref flipFlop425(q[425], d[425], clk, en, clr);
	dffe_ref flipFlop426(q[426], d[426], clk, en, clr);
	dffe_ref flipFlop427(q[427], d[427], clk, en, clr);
	dffe_ref flipFlop428(q[428], d[428], clk, en, clr);
	dffe_ref flipFlop429(q[429], d[429], clk, en, clr);
	dffe_ref flipFlop430(q[430], d[430], clk, en, clr);
	dffe_ref flipFlop431(q[431], d[431], clk, en, clr);
	dffe_ref flipFlop432(q[432], d[432], clk, en, clr);
	dffe_ref flipFlop433(q[433], d[433], clk, en, clr);
	dffe_ref flipFlop434(q[434], d[434], clk, en, clr);
	dffe_ref flipFlop435(q[435], d[435], clk, en, clr);
	dffe_ref flipFlop436(q[436], d[436], clk, en, clr);
	dffe_ref flipFlop437(q[437], d[437], clk, en, clr);
	dffe_ref flipFlop438(q[438], d[438], clk, en, clr);
	dffe_ref flipFlop439(q[439], d[439], clk, en, clr);
	dffe_ref flipFlop440(q[440], d[440], clk, en, clr);
	dffe_ref flipFlop441(q[441], d[441], clk, en, clr);
	dffe_ref flipFlop442(q[442], d[442], clk, en, clr);
	dffe_ref flipFlop443(q[443], d[443], clk, en, clr);
	dffe_ref flipFlop444(q[444], d[444], clk, en, clr);
	dffe_ref flipFlop445(q[445], d[445], clk, en, clr);
	dffe_ref flipFlop446(q[446], d[446], clk, en, clr);
	dffe_ref flipFlop447(q[447], d[447], clk, en, clr);
	dffe_ref flipFlop448(q[448], d[448], clk, en, clr);
	dffe_ref flipFlop449(q[449], d[449], clk, en, clr);
	dffe_ref flipFlop450(q[450], d[450], clk, en, clr);
	dffe_ref flipFlop451(q[451], d[451], clk, en, clr);
	dffe_ref flipFlop452(q[452], d[452], clk, en, clr);
	dffe_ref flipFlop453(q[453], d[453], clk, en, clr);
	dffe_ref flipFlop454(q[454], d[454], clk, en, clr);
	dffe_ref flipFlop455(q[455], d[455], clk, en, clr);
	dffe_ref flipFlop456(q[456], d[456], clk, en, clr);
	dffe_ref flipFlop457(q[457], d[457], clk, en, clr);
	dffe_ref flipFlop458(q[458], d[458], clk, en, clr);
	dffe_ref flipFlop459(q[459], d[459], clk, en, clr);
	dffe_ref flipFlop460(q[460], d[460], clk, en, clr);
	dffe_ref flipFlop461(q[461], d[461], clk, en, clr);
	dffe_ref flipFlop462(q[462], d[462], clk, en, clr);
	dffe_ref flipFlop463(q[463], d[463], clk, en, clr);
	dffe_ref flipFlop464(q[464], d[464], clk, en, clr);
	dffe_ref flipFlop465(q[465], d[465], clk, en, clr);
	dffe_ref flipFlop466(q[466], d[466], clk, en, clr);
	dffe_ref flipFlop467(q[467], d[467], clk, en, clr);
	dffe_ref flipFlop468(q[468], d[468], clk, en, clr);
	dffe_ref flipFlop469(q[469], d[469], clk, en, clr);
	dffe_ref flipFlop470(q[470], d[470], clk, en, clr);
	dffe_ref flipFlop471(q[471], d[471], clk, en, clr);
	dffe_ref flipFlop472(q[472], d[472], clk, en, clr);
	dffe_ref flipFlop473(q[473], d[473], clk, en, clr);
	dffe_ref flipFlop474(q[474], d[474], clk, en, clr);
	dffe_ref flipFlop475(q[475], d[475], clk, en, clr);
	dffe_ref flipFlop476(q[476], d[476], clk, en, clr);
	dffe_ref flipFlop477(q[477], d[477], clk, en, clr);
	dffe_ref flipFlop478(q[478], d[478], clk, en, clr);
	dffe_ref flipFlop479(q[479], d[479], clk, en, clr);
	dffe_ref flipFlop480(q[480], d[480], clk, en, clr);
	dffe_ref flipFlop481(q[481], d[481], clk, en, clr);
	dffe_ref flipFlop482(q[482], d[482], clk, en, clr);
	dffe_ref flipFlop483(q[483], d[483], clk, en, clr);
	dffe_ref flipFlop484(q[484], d[484], clk, en, clr);
	dffe_ref flipFlop485(q[485], d[485], clk, en, clr);
	dffe_ref flipFlop486(q[486], d[486], clk, en, clr);
	dffe_ref flipFlop487(q[487], d[487], clk, en, clr);
	dffe_ref flipFlop488(q[488], d[488], clk, en, clr);
	dffe_ref flipFlop489(q[489], d[489], clk, en, clr);
	dffe_ref flipFlop490(q[490], d[490], clk, en, clr);
	dffe_ref flipFlop491(q[491], d[491], clk, en, clr);
	dffe_ref flipFlop492(q[492], d[492], clk, en, clr);
	dffe_ref flipFlop493(q[493], d[493], clk, en, clr);
	dffe_ref flipFlop494(q[494], d[494], clk, en, clr);
	dffe_ref flipFlop495(q[495], d[495], clk, en, clr);
	dffe_ref flipFlop496(q[496], d[496], clk, en, clr);
	dffe_ref flipFlop497(q[497], d[497], clk, en, clr);
	dffe_ref flipFlop498(q[498], d[498], clk, en, clr);
	dffe_ref flipFlop499(q[499], d[499], clk, en, clr);
	dffe_ref flipFlop500(q[500], d[500], clk, en, clr);
	dffe_ref flipFlop501(q[501], d[501], clk, en, clr);
	dffe_ref flipFlop502(q[502], d[502], clk, en, clr);
	dffe_ref flipFlop503(q[503], d[503], clk, en, clr);
	dffe_ref flipFlop504(q[504], d[504], clk, en, clr);
	dffe_ref flipFlop505(q[505], d[505], clk, en, clr);
	dffe_ref flipFlop506(q[506], d[506], clk, en, clr);
	dffe_ref flipFlop507(q[507], d[507], clk, en, clr);
	dffe_ref flipFlop508(q[508], d[508], clk, en, clr);
	dffe_ref flipFlop509(q[509], d[509], clk, en, clr);
	dffe_ref flipFlop510(q[510], d[510], clk, en, clr);
	dffe_ref flipFlop511(q[511], d[511], clk, en, clr);
	dffe_ref flipFlop512(q[512], d[512], clk, en, clr);
	dffe_ref flipFlop513(q[513], d[513], clk, en, clr);
	dffe_ref flipFlop514(q[514], d[514], clk, en, clr);
	dffe_ref flipFlop515(q[515], d[515], clk, en, clr);
	dffe_ref flipFlop516(q[516], d[516], clk, en, clr);
	dffe_ref flipFlop517(q[517], d[517], clk, en, clr);
	dffe_ref flipFlop518(q[518], d[518], clk, en, clr);
	dffe_ref flipFlop519(q[519], d[519], clk, en, clr);
	dffe_ref flipFlop520(q[520], d[520], clk, en, clr);
	dffe_ref flipFlop521(q[521], d[521], clk, en, clr);
	dffe_ref flipFlop522(q[522], d[522], clk, en, clr);
	dffe_ref flipFlop523(q[523], d[523], clk, en, clr);
	dffe_ref flipFlop524(q[524], d[524], clk, en, clr);
	dffe_ref flipFlop525(q[525], d[525], clk, en, clr);
	dffe_ref flipFlop526(q[526], d[526], clk, en, clr);
	dffe_ref flipFlop527(q[527], d[527], clk, en, clr);
	dffe_ref flipFlop528(q[528], d[528], clk, en, clr);
	dffe_ref flipFlop529(q[529], d[529], clk, en, clr);
	dffe_ref flipFlop530(q[530], d[530], clk, en, clr);
	dffe_ref flipFlop531(q[531], d[531], clk, en, clr);
	dffe_ref flipFlop532(q[532], d[532], clk, en, clr);
	dffe_ref flipFlop533(q[533], d[533], clk, en, clr);
	dffe_ref flipFlop534(q[534], d[534], clk, en, clr);
	dffe_ref flipFlop535(q[535], d[535], clk, en, clr);
	dffe_ref flipFlop536(q[536], d[536], clk, en, clr);
	dffe_ref flipFlop537(q[537], d[537], clk, en, clr);
	dffe_ref flipFlop538(q[538], d[538], clk, en, clr);
	dffe_ref flipFlop539(q[539], d[539], clk, en, clr);
	dffe_ref flipFlop540(q[540], d[540], clk, en, clr);
	dffe_ref flipFlop541(q[541], d[541], clk, en, clr);
	dffe_ref flipFlop542(q[542], d[542], clk, en, clr);
	dffe_ref flipFlop543(q[543], d[543], clk, en, clr);
	dffe_ref flipFlop544(q[544], d[544], clk, en, clr);
	dffe_ref flipFlop545(q[545], d[545], clk, en, clr);
	dffe_ref flipFlop546(q[546], d[546], clk, en, clr);
	dffe_ref flipFlop547(q[547], d[547], clk, en, clr);
	dffe_ref flipFlop548(q[548], d[548], clk, en, clr);
	dffe_ref flipFlop549(q[549], d[549], clk, en, clr);
	dffe_ref flipFlop550(q[550], d[550], clk, en, clr);
	dffe_ref flipFlop551(q[551], d[551], clk, en, clr);
	dffe_ref flipFlop552(q[552], d[552], clk, en, clr);
	dffe_ref flipFlop553(q[553], d[553], clk, en, clr);
	dffe_ref flipFlop554(q[554], d[554], clk, en, clr);
	dffe_ref flipFlop555(q[555], d[555], clk, en, clr);
	dffe_ref flipFlop556(q[556], d[556], clk, en, clr);
	dffe_ref flipFlop557(q[557], d[557], clk, en, clr);
	dffe_ref flipFlop558(q[558], d[558], clk, en, clr);
	dffe_ref flipFlop559(q[559], d[559], clk, en, clr);
	dffe_ref flipFlop560(q[560], d[560], clk, en, clr);
	dffe_ref flipFlop561(q[561], d[561], clk, en, clr);
	dffe_ref flipFlop562(q[562], d[562], clk, en, clr);
	dffe_ref flipFlop563(q[563], d[563], clk, en, clr);
	dffe_ref flipFlop564(q[564], d[564], clk, en, clr);
	dffe_ref flipFlop565(q[565], d[565], clk, en, clr);
	dffe_ref flipFlop566(q[566], d[566], clk, en, clr);
	dffe_ref flipFlop567(q[567], d[567], clk, en, clr);
	dffe_ref flipFlop568(q[568], d[568], clk, en, clr);
	dffe_ref flipFlop569(q[569], d[569], clk, en, clr);
	dffe_ref flipFlop570(q[570], d[570], clk, en, clr);
	dffe_ref flipFlop571(q[571], d[571], clk, en, clr);
	dffe_ref flipFlop572(q[572], d[572], clk, en, clr);
	dffe_ref flipFlop573(q[573], d[573], clk, en, clr);
	dffe_ref flipFlop574(q[574], d[574], clk, en, clr);
	dffe_ref flipFlop575(q[575], d[575], clk, en, clr);
	dffe_ref flipFlop576(q[576], d[576], clk, en, clr);
	dffe_ref flipFlop577(q[577], d[577], clk, en, clr);
	dffe_ref flipFlop578(q[578], d[578], clk, en, clr);
	dffe_ref flipFlop579(q[579], d[579], clk, en, clr);
	dffe_ref flipFlop580(q[580], d[580], clk, en, clr);
	dffe_ref flipFlop581(q[581], d[581], clk, en, clr);
	dffe_ref flipFlop582(q[582], d[582], clk, en, clr);
	dffe_ref flipFlop583(q[583], d[583], clk, en, clr);
	dffe_ref flipFlop584(q[584], d[584], clk, en, clr);
	dffe_ref flipFlop585(q[585], d[585], clk, en, clr);
	dffe_ref flipFlop586(q[586], d[586], clk, en, clr);
	dffe_ref flipFlop587(q[587], d[587], clk, en, clr);
	dffe_ref flipFlop588(q[588], d[588], clk, en, clr);
	dffe_ref flipFlop589(q[589], d[589], clk, en, clr);
	dffe_ref flipFlop590(q[590], d[590], clk, en, clr);
	dffe_ref flipFlop591(q[591], d[591], clk, en, clr);
	dffe_ref flipFlop592(q[592], d[592], clk, en, clr);
	dffe_ref flipFlop593(q[593], d[593], clk, en, clr);
	dffe_ref flipFlop594(q[594], d[594], clk, en, clr);
	dffe_ref flipFlop595(q[595], d[595], clk, en, clr);
	dffe_ref flipFlop596(q[596], d[596], clk, en, clr);
	dffe_ref flipFlop597(q[597], d[597], clk, en, clr);
	dffe_ref flipFlop598(q[598], d[598], clk, en, clr);
	dffe_ref flipFlop599(q[599], d[599], clk, en, clr);
	dffe_ref flipFlop600(q[600], d[600], clk, en, clr);
	dffe_ref flipFlop601(q[601], d[601], clk, en, clr);
	dffe_ref flipFlop602(q[602], d[602], clk, en, clr);
	dffe_ref flipFlop603(q[603], d[603], clk, en, clr);
	dffe_ref flipFlop604(q[604], d[604], clk, en, clr);
	dffe_ref flipFlop605(q[605], d[605], clk, en, clr);
	dffe_ref flipFlop606(q[606], d[606], clk, en, clr);
	dffe_ref flipFlop607(q[607], d[607], clk, en, clr);
	dffe_ref flipFlop608(q[608], d[608], clk, en, clr);
	dffe_ref flipFlop609(q[609], d[609], clk, en, clr);
	dffe_ref flipFlop610(q[610], d[610], clk, en, clr);
	dffe_ref flipFlop611(q[611], d[611], clk, en, clr);
	dffe_ref flipFlop612(q[612], d[612], clk, en, clr);
	dffe_ref flipFlop613(q[613], d[613], clk, en, clr);
	dffe_ref flipFlop614(q[614], d[614], clk, en, clr);
	dffe_ref flipFlop615(q[615], d[615], clk, en, clr);
	dffe_ref flipFlop616(q[616], d[616], clk, en, clr);
	dffe_ref flipFlop617(q[617], d[617], clk, en, clr);
	dffe_ref flipFlop618(q[618], d[618], clk, en, clr);
	dffe_ref flipFlop619(q[619], d[619], clk, en, clr);
	dffe_ref flipFlop620(q[620], d[620], clk, en, clr);
	dffe_ref flipFlop621(q[621], d[621], clk, en, clr);
	dffe_ref flipFlop622(q[622], d[622], clk, en, clr);
	dffe_ref flipFlop623(q[623], d[623], clk, en, clr);
	dffe_ref flipFlop624(q[624], d[624], clk, en, clr);
	dffe_ref flipFlop625(q[625], d[625], clk, en, clr);
	dffe_ref flipFlop626(q[626], d[626], clk, en, clr);
	dffe_ref flipFlop627(q[627], d[627], clk, en, clr);
	dffe_ref flipFlop628(q[628], d[628], clk, en, clr);
	dffe_ref flipFlop629(q[629], d[629], clk, en, clr);
	dffe_ref flipFlop630(q[630], d[630], clk, en, clr);
	dffe_ref flipFlop631(q[631], d[631], clk, en, clr);
	dffe_ref flipFlop632(q[632], d[632], clk, en, clr);
	dffe_ref flipFlop633(q[633], d[633], clk, en, clr);
	dffe_ref flipFlop634(q[634], d[634], clk, en, clr);
	dffe_ref flipFlop635(q[635], d[635], clk, en, clr);
	dffe_ref flipFlop636(q[636], d[636], clk, en, clr);
	dffe_ref flipFlop637(q[637], d[637], clk, en, clr);
	dffe_ref flipFlop638(q[638], d[638], clk, en, clr);
	dffe_ref flipFlop639(q[639], d[639], clk, en, clr);

endmodule