module bitwiseNOT(outR, XR);
	input [31:0] XR;
	output [31:0] outR;

	not a(outR[0], XR[0]);
	not b(outR[1], XR[1]);
	not c(outR[2], XR[2]);
	not d(outR[3], XR[3]);
	not e(outR[4], XR[4]);
	not f(outR[5], XR[5]);
	not g(outR[6], XR[6]);
	not h(outR[7], XR[7]);
	not i(outR[8], XR[8]);
	not j(outR[9], XR[9]);
	not k(outR[10], XR[10]);
	not l(outR[11], XR[11]);
	not m(outR[12], XR[12]);
	not n(outR[13], XR[13]);
	not o(outR[14], XR[14]);
	not p(outR[15], XR[15]);
	not q(outR[16], XR[16]);
	not r(outR[17], XR[17]);
	not s(outR[18], XR[18]);
	not t(outR[19], XR[19]);
	not u(outR[20], XR[20]);
	not v(outR[21], XR[21]);
	not w(outR[22], XR[22]);
	not x(outR[23], XR[23]);
	not y(outR[24], XR[24]);
	not z(outR[25], XR[25]);
	not aa(outR[26], XR[26]);
	not bb(outR[27], XR[27]);
	not cc(outR[28], XR[28]);
	not dd(outR[29], XR[29]);
	not ee(outR[30], XR[30]);
	not ff(outR[31], XR[31]);
	
endmodule