module reg64(q, d, clk, en, clr);
	input [63:0] d; 
	input clk, en, clr;
	output [63:0] q;

	dffe_ref flipFlop0(q[0], d[0], clk, en, clr);
	dffe_ref flipFlop1(q[1], d[1], clk, en, clr);
	dffe_ref flipFlop2(q[2], d[2], clk, en, clr);
	dffe_ref flipFlop3(q[3], d[3], clk, en, clr);
	dffe_ref flipFlop4(q[4], d[4], clk, en, clr);
	dffe_ref flipFlop5(q[5], d[5], clk, en, clr);
	dffe_ref flipFlop6(q[6], d[6], clk, en, clr);
	dffe_ref flipFlop7(q[7], d[7], clk, en, clr);
	dffe_ref flipFlop8(q[8], d[8], clk, en, clr);
	dffe_ref flipFlop9(q[9], d[9], clk, en, clr);
	dffe_ref flipFlop10(q[10], d[10], clk, en, clr);
	dffe_ref flipFlop11(q[11], d[11], clk, en, clr);
	dffe_ref flipFlop12(q[12], d[12], clk, en, clr);
	dffe_ref flipFlop13(q[13], d[13], clk, en, clr);
	dffe_ref flipFlop14(q[14], d[14], clk, en, clr);
	dffe_ref flipFlop15(q[15], d[15], clk, en, clr);
	dffe_ref flipFlop16(q[16], d[16], clk, en, clr);
	dffe_ref flipFlop17(q[17], d[17], clk, en, clr);
	dffe_ref flipFlop18(q[18], d[18], clk, en, clr);
	dffe_ref flipFlop19(q[19], d[19], clk, en, clr);
	dffe_ref flipFlop20(q[20], d[20], clk, en, clr);
	dffe_ref flipFlop21(q[21], d[21], clk, en, clr);
	dffe_ref flipFlop22(q[22], d[22], clk, en, clr);
	dffe_ref flipFlop23(q[23], d[23], clk, en, clr);
	dffe_ref flipFlop24(q[24], d[24], clk, en, clr);
	dffe_ref flipFlop25(q[25], d[25], clk, en, clr);
	dffe_ref flipFlop26(q[26], d[26], clk, en, clr);
	dffe_ref flipFlop27(q[27], d[27], clk, en, clr);
	dffe_ref flipFlop28(q[28], d[28], clk, en, clr);
	dffe_ref flipFlop29(q[29], d[29], clk, en, clr);
	dffe_ref flipFlop30(q[30], d[30], clk, en, clr);
	dffe_ref flipFlop31(q[31], d[31], clk, en, clr);
	dffe_ref flipFlop32(q[32], d[32], clk, en, clr);
	dffe_ref flipFlop33(q[33], d[33], clk, en, clr);
	dffe_ref flipFlop34(q[34], d[34], clk, en, clr);
	dffe_ref flipFlop35(q[35], d[35], clk, en, clr);
	dffe_ref flipFlop36(q[36], d[36], clk, en, clr);
	dffe_ref flipFlop37(q[37], d[37], clk, en, clr);
	dffe_ref flipFlop38(q[38], d[38], clk, en, clr);
	dffe_ref flipFlop39(q[39], d[39], clk, en, clr);
	dffe_ref flipFlop40(q[40], d[40], clk, en, clr);
	dffe_ref flipFlop41(q[41], d[41], clk, en, clr);
	dffe_ref flipFlop42(q[42], d[42], clk, en, clr);
	dffe_ref flipFlop43(q[43], d[43], clk, en, clr);
	dffe_ref flipFlop44(q[44], d[44], clk, en, clr);
	dffe_ref flipFlop45(q[45], d[45], clk, en, clr);
	dffe_ref flipFlop46(q[46], d[46], clk, en, clr);
	dffe_ref flipFlop47(q[47], d[47], clk, en, clr);
	dffe_ref flipFlop48(q[48], d[48], clk, en, clr);
	dffe_ref flipFlop49(q[49], d[49], clk, en, clr);
	dffe_ref flipFlop50(q[50], d[50], clk, en, clr);
	dffe_ref flipFlop51(q[51], d[51], clk, en, clr);
	dffe_ref flipFlop52(q[52], d[52], clk, en, clr);
	dffe_ref flipFlop53(q[53], d[53], clk, en, clr);
	dffe_ref flipFlop54(q[54], d[54], clk, en, clr);
	dffe_ref flipFlop55(q[55], d[55], clk, en, clr);
	dffe_ref flipFlop56(q[56], d[56], clk, en, clr);
	dffe_ref flipFlop57(q[57], d[57], clk, en, clr);
	dffe_ref flipFlop58(q[58], d[58], clk, en, clr);
	dffe_ref flipFlop59(q[59], d[59], clk, en, clr);
	dffe_ref flipFlop60(q[60], d[60], clk, en, clr);
	dffe_ref flipFlop61(q[61], d[61], clk, en, clr);
	dffe_ref flipFlop62(q[62], d[62], clk, en, clr);
	dffe_ref flipFlop63(q[63], d[63], clk, en, clr);

endmodule